../../../IEEE_PROPOSED.src/env_c.vhdl