../../../IEEE_PROPOSED.src/standard_additions_c.vhdl