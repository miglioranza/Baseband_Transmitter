../../../STD.src/standard.vhd