../../../STD.src/textio.vhd