../../../IEEE_PROPOSED.src/standard_textio_additions_c.vhdl